`include "uvm_macros.svh"

package my_env_pkg;
  import uvm_pkg::*;
  import my_agent_pkg::*;
  `include "my_scoreboard.svh"
  `include "my_env.svh"
endpackage : my_env_pkg
